// Prompt: show me a testbench to test the generated bypass fifo bluespec code
// ChatGPT said:
// Here's a Bluespec System Verilog testbench to test your mkBypassFIFO module:

// What this testbench does:
// Enqueues four elements (fills the FIFO).
// Enqueues a fifth element, which should go into bypass.
// Dequeues elements, checking they come out in order.
// Prints values to the console for verification.
                                

package BypassFIFO_Testbench;

import BypassFIFO::*;
import FIFOF::*;
import StmtFSM::*;
import Vector::*;

(* synthesize *)
module mkBypassFIFO_Testbench();

   BypassFIFO#(UInt#(8)) dut <- mkBypassFIFO(UInt#(8), 4);

   Stmt test = 
   seq
      // Enqueue 4 elements
      dut.enq.put(8'h01);
      dut.enq.put(8'h02);
      dut.enq.put(8'h03);
      dut.enq.put(8'h04);

      // Attempt to enqueue 5th element (should trigger bypass)
      dut.enq.put(8'hAA);

      // Dequeue elements
      $display("Dequeue 1: %0h", dut.deq.get);
      dut.deq.deq;
      
      $display("Dequeue 2: %0h", dut.deq.get);
      dut.deq.deq;
      
      $display("Dequeue 3: %0h", dut.deq.get);
      dut.deq.deq;

      $display("Dequeue 4: %0h", dut.deq.get);
      dut.deq.deq;

      // Dequeue bypassed element
      $display("Dequeue Bypassed: %0h", dut.deq.get);
      dut.deq.deq;

      $finish;
   endseq;

   mkAutoFSM(test);

endmodule

endpackage
